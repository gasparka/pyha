library ieee;
    use ieee.fixed_pkg.all;

package ComplexTypes is
end package;
