library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.fixed_float_types.all;
    use ieee.fixed_pkg.all;
    use ieee.math_real.all;

library work;
    use work.all;

package \Register\ is
    type register_t is record
    end record;
    type self_t is record
        \next\: register_t;
    end record;

    procedure reset(reg: inout register_t);
    procedure \__call__\(reg:inout register_t; new_value: unknown_type; ret_0:out unknown_type);
end package;

package body \Register\ is
    procedure reset(reg: inout register_t) is
    begin
    end procedure;

    procedure make_self(reg: register_t; self: out self_t) is
    begin
        self.\next\ := reg;
    end procedure;

    procedure \__call__\(reg:inout register_t; new_value: unknown_type; ret_0:out unknown_type) is
        variable self: self_t;
    begin
        make_self(reg, self);
        self.\next\.a := new_value;
        ret_0 := self.a;
        reg := self.\next\;
    end procedure;
end package body;
