
module top_sv #()
  (
  input clk,rst_n,
  input  [17 :0]    x,
  output [17 :0]    y
  );

  top #()
  top (.*);
endmodule
