library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.fixed_pkg.all;
    use ieee.math_real.all;

library work;
    use work.ComplexTypes.all;
    use work.all;

entity  top is
    port (
        clk, rst_n: in std_logic;

        -- inputs
        in0: in std_logic_vector(37 downto 0);

        -- outputs
        out0: out std_logic_vector(37 downto 0)
    );
end entity;

architecture arch of top is
begin
    process(clk, rst_n)
        variable self: Conjugate_0.register_t;
        -- input variables
        variable var_in0: complex_sfix0_18;

        --output variables
        variable var_out0: complex_sfix0_18;
    begin
    if (not rst_n) then
        Conjugate_0.reset(self);
    elsif rising_edge(clk) then
        --convert slv to normal types
        var_in0 := (real=>to_sfixed(in0(37 downto 19), 0, -18), imag=>to_sfixed(in0(18 downto 0), 0, -18));

        --call the main entry
        Conjugate_0.main(self, var_in0, ret_0=>var_out0);

        --convert normal types to slv
        out0 <= to_slv(var_out0.real) & to_slv(var_out0.imag);
      end if;

    end process;
end architecture;