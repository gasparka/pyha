--library ieee;
--  use ieee.std_logic_1164.all;
--  use ieee.numeric_std.all;
--  use ieee.numeric_std.all;
--  use ieee.fixed_float_types.all;
--  use ieee.fixed_pkg.all;

--package PyhaUtil is
--  type sfixed_list_t is array (natural range <>) of sfixed;
-- type integer_list_t is array (natural range <>) of integer;
--  type boolean_list_t is array (natural range <>) of boolean;
--end package;

package Util is
  type integer_list_t is array (natural range <>) of integer;
end package;