
module top_sv #()
  (
  input clk,rst_n,
  input  [27 :0]    in0,
  output [27 :0]    out0
  );

  top #()
  top (.*);
endmodule
