
module top_sv #()
  (
  input clk,rst_n,
  input  [17 :0]    x1,
  output [17 :0]    y1
  );

  top #()
  top (.*);
endmodule
