
module top_sv #()
  (
  input clk,rst_n,
  input  [17 :0]    x1,x2,
  output [17 :0]    y1,y2
  );

  top #()
  top (.*);
endmodule
